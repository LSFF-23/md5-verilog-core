module fmax_wiring (clk, rst_n, start, sel, out, done);
input clk, rst_n, start;
input sel;
output [0:127] out;
output done;

reg [0:511] s512 [1:0];
wire core_resume;

assign core_resume = start & done ;

md5_core core (clk, rst_n, start, core_resume, s512[sel], out, done);

initial begin
    s512[0] = 512'h58585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858;
    s512[1] = 512'h58585858585858585858585858585858585858585858585858585858585858585858585880000000000000000000000000000000000000002003000000000000;
end

endmodule