module tb_md5_core;
reg clk, h_rst, s_rst;
reg [0:511] input_data;
wire [0:127] hash;
wire done;

md5_core dut (clk, h_rst, s_rst, input_data, hash, done);

always #5 clk = !clk;

initial begin
    clk = 0; h_rst = 0; s_rst = 0; #10

    input_data = 512'h58585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858585858;
    h_rst = 1; #10
    h_rst = 0; #690

    input_data = 512'h58585858585858585858585858585858585858585858585858585858585858585858585880000000000000000000000000000000000000002003000000000000;
    s_rst = 1; #10
    s_rst = 0; #690
    $stop(0);
end

endmodule